`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "mem_common.sv"
`include "mem_tx.sv"

`include "mem_sequencer.sv"
`include "mem_driver.sv"
`include "mem_monitor.sv"
`include "mem_coverage.sv"

`include "mem_sbd.sv"
`include "mem_agent.sv"
`include "mem_env.sv"

`include "test_lib.sv"
`include "top.sv"

